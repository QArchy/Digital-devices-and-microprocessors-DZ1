library verilog;
use verilog.vl_types.all;
entity count_down_vlg_vec_tst is
end count_down_vlg_vec_tst;
