library verilog;
use verilog.vl_types.all;
entity a_chema is
    port(
        y_a             : out    vl_logic;
        x3              : in     vl_logic;
        x2              : in     vl_logic;
        x0              : in     vl_logic;
        x1              : in     vl_logic
    );
end a_chema;
