library verilog;
use verilog.vl_types.all;
entity g_schema_vlg_vec_tst is
end g_schema_vlg_vec_tst;
