library verilog;
use verilog.vl_types.all;
entity y_a_vlg_vec_tst is
end y_a_vlg_vec_tst;
