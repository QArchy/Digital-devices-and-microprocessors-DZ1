library verilog;
use verilog.vl_types.all;
entity a_chema_vlg_check_tst is
    port(
        y_a             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end a_chema_vlg_check_tst;
