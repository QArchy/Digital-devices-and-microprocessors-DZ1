library verilog;
use verilog.vl_types.all;
entity CNT_without_R_vlg_vec_tst is
end CNT_without_R_vlg_vec_tst;
