library verilog;
use verilog.vl_types.all;
entity d_schema_vlg_vec_tst is
end d_schema_vlg_vec_tst;
