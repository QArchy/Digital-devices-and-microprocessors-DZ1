library verilog;
use verilog.vl_types.all;
entity BCD_after_CNT_vlg_vec_tst is
end BCD_after_CNT_vlg_vec_tst;
