library verilog;
use verilog.vl_types.all;
entity c_schema_vlg_vec_tst is
end c_schema_vlg_vec_tst;
