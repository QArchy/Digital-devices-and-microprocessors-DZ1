library verilog;
use verilog.vl_types.all;
entity b_schema is
    port(
        b               : out    vl_logic;
        x3              : in     vl_logic;
        x2              : in     vl_logic;
        x0              : in     vl_logic;
        x1              : in     vl_logic
    );
end b_schema;
