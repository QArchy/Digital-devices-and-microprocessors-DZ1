library verilog;
use verilog.vl_types.all;
entity c_schema_vlg_check_tst is
    port(
        y_c             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end c_schema_vlg_check_tst;
