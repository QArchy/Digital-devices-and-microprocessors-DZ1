library verilog;
use verilog.vl_types.all;
entity Counter_to_6_vlg_vec_tst is
end Counter_to_6_vlg_vec_tst;
