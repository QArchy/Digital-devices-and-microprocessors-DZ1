library verilog;
use verilog.vl_types.all;
entity e_schema_vlg_vec_tst is
end e_schema_vlg_vec_tst;
