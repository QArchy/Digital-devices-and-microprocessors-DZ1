library verilog;
use verilog.vl_types.all;
entity f_schema_vlg_vec_tst is
end f_schema_vlg_vec_tst;
