library verilog;
use verilog.vl_types.all;
entity f_schema_vlg_check_tst is
    port(
        y_f             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end f_schema_vlg_check_tst;
