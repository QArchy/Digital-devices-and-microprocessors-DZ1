library verilog;
use verilog.vl_types.all;
entity Frequency_divider_vlg_vec_tst is
end Frequency_divider_vlg_vec_tst;
