library verilog;
use verilog.vl_types.all;
entity b_schema_vlg_vec_tst is
end b_schema_vlg_vec_tst;
