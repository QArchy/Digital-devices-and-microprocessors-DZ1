library verilog;
use verilog.vl_types.all;
entity Counter_to_6_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Counter_to_6_vlg_sample_tst;
