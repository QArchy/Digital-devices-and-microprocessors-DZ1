library verilog;
use verilog.vl_types.all;
entity test3 is
    port(
        Q0              : out    vl_logic;
        c               : in     vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic
    );
end test3;
