library verilog;
use verilog.vl_types.all;
entity test2_vlg_sample_tst is
    port(
        c               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end test2_vlg_sample_tst;
