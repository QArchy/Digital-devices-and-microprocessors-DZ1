library verilog;
use verilog.vl_types.all;
entity Freq_divider_vlg_vec_tst is
end Freq_divider_vlg_vec_tst;
