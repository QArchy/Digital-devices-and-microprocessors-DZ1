library verilog;
use verilog.vl_types.all;
entity test_sub_vlg_check_tst is
    port(
        pin_name2       : in     vl_logic;
        pin_name3       : in     vl_logic;
        pin_name4       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end test_sub_vlg_check_tst;
