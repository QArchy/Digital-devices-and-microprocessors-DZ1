library verilog;
use verilog.vl_types.all;
entity test3_vlg_sample_tst is
    port(
        c               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end test3_vlg_sample_tst;
