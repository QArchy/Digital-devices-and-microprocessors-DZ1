library verilog;
use verilog.vl_types.all;
entity recoder_schema_vlg_vec_tst is
end recoder_schema_vlg_vec_tst;
