library verilog;
use verilog.vl_types.all;
entity count_down_vlg_check_tst is
    port(
        y0              : in     vl_logic;
        y1              : in     vl_logic;
        y2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end count_down_vlg_check_tst;
