library verilog;
use verilog.vl_types.all;
entity recoder_schema_vlg_sample_tst is
    port(
        Q0              : in     vl_logic;
        Q1              : in     vl_logic;
        Q2              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end recoder_schema_vlg_sample_tst;
