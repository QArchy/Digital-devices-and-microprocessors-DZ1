library verilog;
use verilog.vl_types.all;
entity d_schema_vlg_check_tst is
    port(
        y_d             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end d_schema_vlg_check_tst;
