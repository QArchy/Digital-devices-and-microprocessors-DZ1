library verilog;
use verilog.vl_types.all;
entity e_schema is
    port(
        y_e             : out    vl_logic;
        x3              : in     vl_logic;
        x1              : in     vl_logic;
        x0              : in     vl_logic;
        x2              : in     vl_logic
    );
end e_schema;
