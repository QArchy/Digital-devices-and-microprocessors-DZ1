library verilog;
use verilog.vl_types.all;
entity counter3Bit_reset_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end counter3Bit_reset_vlg_sample_tst;
