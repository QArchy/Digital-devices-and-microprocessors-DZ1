library verilog;
use verilog.vl_types.all;
entity counter3Bit_reset_vlg_vec_tst is
end counter3Bit_reset_vlg_vec_tst;
