library verilog;
use verilog.vl_types.all;
entity test2 is
    port(
        pin_name2       : out    vl_logic;
        c               : in     vl_logic
    );
end test2;
