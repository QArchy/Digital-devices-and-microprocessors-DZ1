library verilog;
use verilog.vl_types.all;
entity g_schema_vlg_check_tst is
    port(
        y_g             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g_schema_vlg_check_tst;
