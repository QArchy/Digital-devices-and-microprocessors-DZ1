library verilog;
use verilog.vl_types.all;
entity e_schema_vlg_check_tst is
    port(
        y_e             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end e_schema_vlg_check_tst;
