library verilog;
use verilog.vl_types.all;
entity c_schema is
    port(
        y_c             : out    vl_logic;
        x3              : in     vl_logic;
        x2              : in     vl_logic;
        x0              : in     vl_logic;
        x1              : in     vl_logic
    );
end c_schema;
