library verilog;
use verilog.vl_types.all;
entity BCD_schema_vlg_vec_tst is
end BCD_schema_vlg_vec_tst;
