library verilog;
use verilog.vl_types.all;
entity CNT1_vlg_vec_tst is
end CNT1_vlg_vec_tst;
