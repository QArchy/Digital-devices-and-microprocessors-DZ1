library verilog;
use verilog.vl_types.all;
entity CNT_v_vlg_vec_tst is
end CNT_v_vlg_vec_tst;
