library verilog;
use verilog.vl_types.all;
entity Test2_vlg_sample_tst is
    port(
        C               : in     vl_logic;
        PRN             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Test2_vlg_sample_tst;
