library verilog;
use verilog.vl_types.all;
entity c_schema_vlg_sample_tst is
    port(
        x0              : in     vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end c_schema_vlg_sample_tst;
