library verilog;
use verilog.vl_types.all;
entity a_chema_vlg_vec_tst is
end a_chema_vlg_vec_tst;
