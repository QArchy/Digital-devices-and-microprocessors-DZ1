library verilog;
use verilog.vl_types.all;
entity RS_vlg_vec_tst is
end RS_vlg_vec_tst;
