library verilog;
use verilog.vl_types.all;
entity counter5Bit_verilog_schema_vlg_vec_tst is
end counter5Bit_verilog_schema_vlg_vec_tst;
