library verilog;
use verilog.vl_types.all;
entity counter5Bit_verilog_schema_vlg_check_tst is
    port(
        Q_1             : in     vl_logic;
        Q_2             : in     vl_logic;
        Q_3             : in     vl_logic;
        Q_4             : in     vl_logic;
        Q_5             : in     vl_logic;
        Q_6             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end counter5Bit_verilog_schema_vlg_check_tst;
