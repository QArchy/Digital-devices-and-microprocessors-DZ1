library verilog;
use verilog.vl_types.all;
entity Test2_vlg_vec_tst is
end Test2_vlg_vec_tst;
